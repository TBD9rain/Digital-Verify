//==================================================================================================
//
//  Project         :   Digital Verify Example
//  Version         :   v1.0.0
//  Title           :   verify_pkg
//
//  Description     :   package components for Verification
//
//  Additional info :
//  Author          :   lshi1
//  Email           :
//
//==================================================================================================

package verify_pkg;

import msg_log_pkg::*;

//  specify the relative path from simulation work directory
`include "../sim/../tb/test_ifc.sv"
`include "../sim/../tb/test_cls.sv"


endpackage

